package packet_pkg;

 // `include "port_if.sv"  
   // `include "switch_port.sv" 
 `include "packet_data.sv"
  
  `include "component_base.sv"

 
  `include "sequencer.sv" 
  `include "driver.sv"      
  `include "monitor.sv"     

  `include "agent.sv"      
  `include "packet_vc.sv"  

endpackage

